//Project: RISC-V 32 bit Architecture
//Module: tb_Program_Counter (FU)
//Author: Sistla Manojna
//Updated: 06/03/2020
//Updates the Program Counter value
//Updates:

module tb_Program_Counter();
endmodule
